module fifo_sync (
    input logic clk,
    input logic rd,
    input logic wr,
    
    output logic full,
    output logic empty
);
    

always @(posedge clk) begin
    
end

endmodule